---------------------------------------------------------
--									PLDP
--								  A N E M
--
--						Test Bench do banco de registradores
--
--					Bruno Morais / Lucas Lessa
---------------------------------------------------------
--Utiliza entidade externa BancoReg (Banco de registradores)
-- : BancoReg.vhd			
---------------------------------------------------------

--Data ult. mod.	:	02/05/2011
--Changelog:
---------------------------------------------------------
--@02/05/2011: Versão inicial

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;

ENTITY REG_FILE_TB IS

--GENERICOS PARA CONFIGURAR O TAMANHO DOS DADOS DOS REGISTRADORES E TAMANHO DO BANCO
GENERIC( N: NATURAL := 16; P: NATURAL := 8; Q: NATURAL := 4);

END REG_FILE_TB;

ARCHITECTURE BEHAVIOR OF REG_FILE_TB IS

--SINAIS INTERNOS PARA CONEXAO COM O BANCO DE REGISTRADORES
SIGNAL S_IN,TEST,CK,RST,S_OUT: STD_LOGIC := '0';
SIGNAL ULA_IN,DATA_IN,A_OUT,B_OUT: STD_LOGIC_VECTOR( N-1 DOWNTO 0) := (OTHERS=>'0');
SIGNAL BYTE_IN: STD_LOGIC_VECTOR(P-1 DOWNTO 0) := (OTHERS=>'0');
SIGNAL SEL_A,SEL_B: STD_LOGIC_VECTOR(Q-1 DOWNTO 0) := "0000";
SIGNAL REG_CNT: STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
  

BEGIN

--BANCO DE REGISTRADORES
  
REGBNK : ENTITY WORK.BANCOREG(ANEM) GENERIC MAP(W=>P,DATA_W=>N,REGBNK_ADDR=>Q,REGBNK_SIZE=>N) 
  PORT MAP(S_IN=>S_IN,TEST=>TEST,ULA_IN=>ULA_IN,BYTE_IN=>BYTE_IN,SEL_A=>SEL_A,SEL_B=>SEL_B,DATA_IN=>DATA_IN,CK=>CK,RST=>RST,REG_CNT=>REG_CNT,A_OUT=>A_OUT,B_OUT=>B_OUT,S_OUT=>S_OUT);
  
PROCESS
    
--PREPARA PARA CARREGAR ARQUIVO COM DADOS DE TESTE
FILE ARQUIVO: TEXT IS IN "teste.prn";

VARIABLE    LINHA: LINE; --UMA LINHA DO ARQUIVO
VARIABLE ENDERECO: BIT_VECTOR(3 DOWNTO 0) := (OTHERS=>'0'); --ENDERECO DO REGISTRADOR NO BANCO
VARIABLE    DADOS: BIT_VECTOR(15 DOWNTO 0) := (OTHERS=>'0'); --DADOS
VARIABLE      SEL: BIT_VECTOR(2 DOWNTO 0) := (OTHERS=>'0'); --CONTROLE DE OPERACOES

--SINAIS NAO RECEBEM IMEDIATAMENTE SEUS VALORES!
    
BEGIN
  
  --RESETA BANCO DE REGISTRADORES MANUALMENTE
  
    RST <= '1';
  
    WAIT FOR 10ns;
  
    RST<= '0';
  
    WAIT FOR 10ns;
    
  --LOOP DE LEITURA E TESTES
  
  WHILE (NOT ENDFILE(ARQUIVO)) LOOP
    

	--REALIZA LEITURA E  TESTES QUANDO O CLOCK ESTA ALTO, PARA COMPENSAR
	--O ATRASO DE RECEBIMENTO DOS SINAIS
	
	--SO TESTA REG_A, POIS OS DADOS SAO GRAVADOS APENAS NELE.
    
  IF CK = '1' THEN 
    
    --LE UMA LINHA
    
    READLINE(ARQUIVO,LINHA);
    
    --LE DADOS DA LINHA
    
    READ(LINHA,ENDERECO);
    READ(LINHA,DADOS);
    READ(LINHA,SEL);
    
    --COLOCA O ENDERECO LIDO DA LINHA EM SEL_A
    --NOTA: O SINAL SEL_A SO TEM O VALOR "ENDERECO" NO PROXIMO CICLO!
    
    SEL_A   <= TO_STDLOGICVECTOR(ENDERECO);
    
    --COLOCA OS BITS DE CONTROLE EM REG_CNT
    
    REG_CNT <= TO_STDLOGICVECTOR(SEL);
    
    --COLOCA OS DADOS LIDOS TANTO EM DATA_IN QUANTO EM ULA_IN,
    --QUEM VAI DECIDIR QUAL DOS DOIS SERA UTILIZADO E O BANCO,
    --DEPENDENDO DE REG_CNT

    DATA_IN <= TO_STDLOGICVECTOR(DADOS);
    ULA_IN <= TO_STDLOGICVECTOR(DADOS);
    
    --VERIFICA SE ESTA COLOCANDO UM VALOR BYTE A BYTE
    
    IF SEL = "010" THEN
    
		--COLOCANDO VALOR NO BYTE SUPERIOR DE REG_A
      
        BYTE_IN <= TO_STDLOGICVECTOR(DADOS)(15 DOWNTO 8);
      
    ELSIF SEL = "011" THEN
    
		--COLOCANDO VALOR NO BYTE INFERIOR DE REG_B
    
        BYTE_IN <= TO_STDLOGICVECTOR(DADOS)(7 DOWNTO 0);
      
    ELSE BYTE_IN <= (OTHERS=>'0'); --ZERA BYTE_IN, EVITA LATCHES
    
 END IF;  
 
 END IF;  
 
  --CLOCK

  WAIT FOR 10NS;
  
  CK <= NOT CK;
  
END LOOP;

  --MAIS UM CLOCK PARA REGISTRAR O ULTIMO VALOR COLOCADO

  WAIT FOR 10NS;
  
  CK <= NOT CK;
    
END PROCESS;

END ARCHITECTURE;
   


