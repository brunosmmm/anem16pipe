LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE STD.TEXTIO.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Debug IS

    GENERIC (INST_END_SIZE : INTEGER := 16;
             MSG_MAX_SIZE : INTEGER := 32);
    
    PORT ( INST_END : STD_LOGIC_VECTOR(INST_END_SIZE-1 DOWNTO 0));
           
END ENTITY;

ARCHITECTURE ANEM OF Debug IS

TYPE DEBUG_MSGS IS ARRAY(((2**INST_END_SIZE)-1) DOWNTO 0) OF STRING(1 TO MSG_MAX_SIZE);
SIGNAL MESSAGES : DEBUG_MSGS;

BEGIN

MAIN: PROCESS

    FILE DEBUGMSG : TEXT IS IN "debug.txt";
    VARIABLE LINHA: LINE;
    VARIABLE ADDR : BIT_VECTOR(INST_END_SIZE-1 DOWNTO 0);
    VARIABLE MSG : STRING(1 TO MSG_MAX_SIZE);
    
    BEGIN
    
        WHILE NOT ENDFILE(DEBUGMSG) LOOP
        
            READLINE(DEBUGMSG,LINHA);
            READ(LINHA,ADDR);

            READ(LINHA,MSG);
            
            MESSAGES(conv_integer(to_stdlogicvector(ADDR))) <= MSG; 
            
        END LOOP;
        
END PROCESS;
    
DBG: PROCESS(INST_END) 
    
    BEGIN
     
    IF MESSAGES(conv_integer(INST_END)) /= "0000000000000000000000000000000" THEN
    
        REPORT(MESSAGES(conv_integer(INST_END)));
        
    END IF;
       
END PROCESS;

END ARCHITECTURE;
