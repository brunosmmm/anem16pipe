-----------------------------
--! @file test_bench.vhd
--! @brief ANEM test bench
--! @date 2011,2014
-----------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TEST_BENCH IS
  GENERIC( N: NATURAL := 256);
END TEST_BENCH;

ARCHITECTURE TESTE OF TEST_BENCH IS

  SIGNAL CK, RST: STD_LOGIC := '0';
  SIGNAL INST: STD_LOGIC_VECTOR(15 DOWNTO 0);  --! next instruction
  SIGNAL INST_ADDR: STD_LOGIC_VECTOR(15 DOWNTO 0):= (OTHERS => '0'); --! next instruction address
  SIGNAL TEST: STD_LOGIC := '0';  --! test mode enable
  SIGNAL MEM_W: STD_LOGIC;     --! memory write enable
  SIGNAL MEM_EN: STD_LOGIC;    --! memory enable

  SIGNAL DATA : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS=>'Z'); --! bidirectional data bus

  SIGNAL MEM_ADDR: STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL BIT_INST_OUT: STD_LOGIC;

  -- GPIO pins
  signal porta_pins : std_logic_vector(15 downto 0) := (others => 'Z');
  signal portb_pins : std_logic_vector(15 downto 0) := (others => 'Z');

BEGIN

  cpu:  entity work.ANEM(test)
    PORT MAP(CK=>CK,
             RST=>RST,
             TEST=>TEST,
             INST=>INST,
             S_IN=>'0',
             S_OUT=>BIT_INST_OUT,
             MEM_W=>MEM_W,
             MEM_EN=>MEM_EN,
             MEM_ADDR=>MEM_ADDR,
             DATA=>DATA,
             INST_ADDR=>INST_ADDR,
             INT=>'0'
             );

  imem: entity work.progmem(rom)
    PORT MAP(ck=>CK,
             en=>'1',
             address=>INST_ADDR,
             instr=>INST
             );

  dmem: entity work.datamem(ram)
    PORT MAP(ck=>CK,
             en=>MEM_EN,
             w=>MEM_W,
             address=>MEM_ADDR,
             data=>DATA);

  -- MAC peripheral
  mac_inst: ENTITY WORK.MAC(MultAcc)
    PORT MAP(DATA=>DATA, CK=>CK, RST=>RST, ADDR=>MEM_ADDR,
             W=>MEM_W, EN=>MEM_EN, INT=>OPEN);

  -- GPIO peripheral
  gpio_inst: entity work.gpio(behavioral)
    port map(DATA=>DATA, ADDR=>MEM_ADDR, W=>MEM_W, EN=>MEM_EN,
             CK=>CK, RST=>RST, PORTA_PINS=>porta_pins,
             PORTB_PINS=>portb_pins, INT=>open);

  -- Timer peripheral
  timer_inst: entity work.timer(behavioral)
    port map(DATA=>DATA, ADDR=>MEM_ADDR, W=>MEM_W, EN=>MEM_EN,
             CK=>CK, RST=>RST, INT=>open);

  -- UART peripheral
  uart_inst: entity work.uart(behavioral)
    port map(DATA=>DATA, ADDR=>MEM_ADDR, W=>MEM_W, EN=>MEM_EN,
             CK=>CK, RST=>RST, TX=>open, RX=>'1', INT=>open);

  PROCESS

  begin

    RST <=  '1';
    WAIT FOR 30NS;
    RST <=  '0';

    FOR I IN 0 TO 2048 LOOP                -- clk
      CK <= NOT CK;
      WAIT FOR 10 NS;
    END LOOP;
  END PROCESS;
END TESTE;
